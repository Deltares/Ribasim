netcdf basin_state {
dimensions:
	time = 1 ;
	stations = 6 ;
	char_leng_id = 64 ;
	char_leng_name = 255 ;
variables:
	double time(time) ;
		string time:standard_name = "time" ;
		string time:long_name = "time" ;
		string time:units = "minutes since 1970-01-01 00:00:00.0 +0000" ;
		string time:axis = "T" ;
	double lat(stations) ;
		string lat:standard_name = "latitude" ;
		string lat:long_name = "Station coordinates, latitude" ;
		string lat:units = "degrees_north" ;
		string lat:axis = "Y" ;
		lat:_FillValue = 9.96921e+036 ;
	double lon(stations) ;
		string lon:standard_name = "longitude" ;
		string lon:long_name = "Station coordinates, longitude" ;
		string lon:units = "degrees_east" ;
		string lon:axis = "X" ;
		lon:_FillValue = 9.96921e+036 ;
	double y(stations) ;
		string y:standard_name = "latitude" ;
		string y:long_name = "y coordinate according to WGS 1984" ;
		string y:units = "degrees_north" ;
		string y:axis = "Y" ;
		y:_FillValue = 9.96921e+036 ;
	double x(stations) ;
		string x:standard_name = "longitude" ;
		string x:long_name = "x coordinate according to WGS 1984" ;
		string x:units = "degrees_east" ;
		string x:axis = "X" ;
		x:_FillValue = 9.96921e+036 ;
	double z(stations) ;
		string z:long_name = "height above mean sea level" ;
		string z:units = "meters" ;
		z:_FillValue = 9.96921e+036 ;
	char station_id(stations, char_leng_id) ;
		string station_id:long_name = "station identification code" ;
		string station_id:cf_role = "timeseries_id" ;
	char station_names(stations, char_leng_name) ;
		string station_names:long_name = "station name" ;
	float level(time, stations) ;
		string level:long_name = "level" ;
		string level:units = "m" ;
		level:_FillValue = -999.f ;
		string level:coordinates = "lat lon x y z station_id" ;

// global attributes:
		string :Conventions = "CF-1.6" ;
		string :title = "Data" ;
		string :institution = "Deltares" ;
		string :source = "Export NETCDF-CF_TIMESERIES from Delft-FEWS" ;
		string :history = "2026-01-14 09:36:58 GMT: exported from Delft-FEWS" ;
		string :references = "http://www.delft-fews.com" ;
		string :Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		string :summary = "Data exported from Delft-FEWS" ;
		string :date_created = "2026-01-14 09:36:58 GMT" ;
		string :fews_implementation_version = "2025.01" ;
		string :fews_patch_number = "509261311" ;
		string :fews_build_number = "508210944" ;
		string :coordinate_system = "WGS 1984" ;
		string :featureType = "timeSeries" ;
		string :time_coverage_start = "2025-11-05T00:00:00+0000" ;
		string :time_coverage_end = "2025-11-05T00:00:00+0000" ;
		string :geospatial_lon_min = "99.068673" ;
		string :geospatial_lon_max = "99.643538" ;
		string :geospatial_lat_min = "17.499098" ;
		string :geospatial_lat_max = "18.809239" ;
data:

 time = 29371680 ;

 lat = 52.0, 52.1, 52.2, 52.3, 52.4, 52.5 ;

 lon = 5.1, 5.2, 5.3, 5.4, 5.5, 5.6 ;

 y = 52.0, 52.1, 52.2, 52.3, 52.4, 52.5 ;

 x = 5.1, 5.2, 5.3, 5.4, 5.5, 5.6 ;

 z = 0, 0, 0, 0, 0, 0 ;

 station_id =
  "101",
  "102",
  "103",
  "104",
  "105",
  "106" ;

 station_names =
  "basin_a",
  "basin_b",
  "basin_c",
  "basin_d",
  "basin_e",
  "basin_f" ;

 level =
  1.1, 1.2, 1.3, 1.4, 1.5, 1.6 ;
}
